module my_not(
    input a,
    output y
  );
  assign y=~a;
endmodule

